SoC_Map.bsv